`timescale 1ns / 1ps // <simulation time step> / <simulation time step precision>
//////////////////////////////////////////////////////////////////////////////////
// Firmware to drive a MAX5875 DAC in interleaved mode
//
// Daniel Schussheim
//////////////////////////////////////////////////////////////////////////////////
module MAX5875(
    input wire clk_in,
    input wire signed [15:0] s_in0,
    input wire signed [15:0] s_in1,
    output wire clk_out,
    output reg sel,
    output reg signed [15:0] s_out
);
// Output clock to DACs
assign clk_out = clk_in;

// sel and sel_int are (100 MHz) channel selects. Because sel is an output to the DAC, implementation forces it to be generated by a flip-flop (FF) in an I/O Block (IOB), whereas sel_int has to be generated by a fabric FF to be used internally in the FPGA.
// This avoids using a FF in an IOB to drive signals in the logical fabric or other IOB's, which causes a placement error.
// Including a DONT_TOUCH synthesis directive before the below declaration of sel_int prevents the optimization of sel and sel_int into a single signal before placement.
(* DONT_TOUCH = "TRUE" *)
reg sel_int = 1'b0;
// "DDR" data output (update in between sel changes)
always @(posedge clk_in) begin
sel_int <= !sel_int;
sel     <= !sel_int;
    if (sel_int)
        s_out <= s_in1;
    else
        s_out <= s_in0;
end

endmodule
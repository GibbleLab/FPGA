    phs0 = 33.75,   phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 213.75,  phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 264.375, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 354.375, phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 292.5,   phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 56.25,   phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 39.375,  phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 315,     phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 241.875, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 11.25,   phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 264.375, phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 286.875, phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 168.75,  phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 298.125, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 135,     phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 118.125, phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 264.375, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 0,       phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 5.625,   phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 343.125, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 326.25,  phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 129.375, phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 5.625,   phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 90,      phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 315,     phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 90,      phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 225,     phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 253.125, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 84.375,  phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 253.125, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 33.75,   phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 61.875,  phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 56.25,   phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 174.375, phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 140.625, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 303.75,  phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 135,     phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 140.625, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 303.75,  phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 326.25,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 28.125,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 112.5,   phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 281.25,  phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 84.375,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 135,     phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 174.375, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 241.875, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 11.25,   phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 258.75,  phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 298.125, phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 157.5,   phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 354.375, phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 219.375, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 241.875, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 123.75,  phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 174.375, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 157.5,   phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 247.5,   phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 281.25,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 309.375, phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 50.625,  phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 168.75,  phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 281.25,  phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 354.375, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 286.875, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 118.125, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 163.125, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 286.875, phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 174.375, phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 163.125, phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 253.125, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 129.375, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 0,       phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 219.375, phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 78.75,   phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 343.125, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 281.25,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 151.875, phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 146.25,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 151.875, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 331.875, phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 354.375, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 264.375, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 101.25,  phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 315,     phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 286.875, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 61.875,  phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 258.75,  phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 185.625, phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 67.5,    phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 241.875, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 202.5,   phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 303.75,  phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 140.625, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 123.75,  phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 90,      phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 123.75,  phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 258.75,  phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 90,      phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 208.125, phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 0,     phs5 = 0, phs6 = 123.75;
    phs0 = 337.5,   phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 196.875, phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 331.875, phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 129.375, phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 253.125, phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 84.375,  phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 101.25,  phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 208.125, phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 67.5,    phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 281.25,  phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 28.125,  phs1 = 0, phs2 = 0, phs3 = 22.5,  phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 56.25,   phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 157.5, phs5 = 0, phs6 = 123.75;
    phs0 = 303.75,  phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 315,     phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 337.5,   phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 202.5,   phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 151.875, phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 22.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 253.125, phs1 = 0, phs2 = 0, phs3 = 90,    phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 298.125, phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 16.875,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 281.25,  phs1 = 0, phs2 = 0, phs3 = 45,    phs4 = 45,    phs5 = 0, phs6 = 123.75;
    phs0 = 11.25,   phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 213.75,  phs1 = 0, phs2 = 0, phs3 = 112.5, phs4 = 135,   phs5 = 0, phs6 = 123.75;
    phs0 = 28.125,  phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 90,    phs5 = 0, phs6 = 123.75;
    phs0 = 33.75,   phs1 = 0, phs2 = 0, phs3 = 157.5, phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 174.375, phs1 = 0, phs2 = 0, phs3 = 135,   phs4 = 112.5, phs5 = 0, phs6 = 123.75;
    phs0 = 196.875, phs1 = 0, phs2 = 0, phs3 = 0,     phs4 = 67.5,  phs5 = 0, phs6 = 123.75;
    phs0 = 95.625,  phs1 = 0, phs2 = 0, phs3 = 67.5,  phs4 = 135,   phs5 = 0, phs6 = 123.75;
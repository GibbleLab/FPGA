    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 1, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 1, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 1, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 1, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 1; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 3, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 3, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 3, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 3, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 3; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 5, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 5, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 5, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 5, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 5; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 7, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 7, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 7, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 7, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 7; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 9, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 9, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 9, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 9, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 9; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 11, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 11, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 11, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 11, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 11; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 13, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 13, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 13, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 13, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 13; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 15, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 15, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 15, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 15, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 15; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 17, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 17, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 17, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 17, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 17; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 19, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 19, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 19, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 19, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 19; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 21, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 21, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 21, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 21, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 21; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 23, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 23, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 23, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 23, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 23; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 25, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 25, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 25, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 25, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 25; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 27, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 27, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 27, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 27, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 27; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 29, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 29, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 29, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 29, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 29; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])

    dly00 = 8,  dly01 = 9,  dly10 = 10, dly11 = 9,  dlyf0 = 31, // delays for D00[0], D00[1], D01[0], D01[1], FR0 ([,], [,], [,], [,], [,])
    dly20 = 22, dly21 = 23, dly30 = 24, dly31 = 24, dlyf1 = 31, // delays for D10[0], D10[1], D11[0], D11[1], FR1 ([,], [,], [,], [,], [,])
    dly40 = 19, dly41 = 15, dly50 = 14, dly51 = 13, dlyf2 = 31, // delays for D20[0], D20[1], D21[0], D21[1], FR2 ([,], [,], [,], [,], [,])
    dly60 = 14, dly61 = 16, dly70 = 17, dly71 = 17, dlyf3 = 31, // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
    dly80 = 16, dly81 = 17, dly90 = 16, dly91 = 16, dlyf4 = 31; // delays for D30[0], D30[1], D31[0], D31[1], FR3 ([,], [,], [,], [,], [,])
